module PC_REG(
    input logic clk,
    input logic rst,
    input logic [31:0] next_PC,
    output logic [31:0] PC
);



endmodule

