module ALU(
    input logic [31:0] ALU_Op1,
    input logic [31:0] ALU_Op2,
    input logic [2:0] ALUctrl,
    output logic [31:0] ALU_out,
    output logic EQ
);



endmodule


