module InstrMem(
    input logic [31:0] Imem_Addr,
    output logic [31:0] Read_Data
);



endmodule

