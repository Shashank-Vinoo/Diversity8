module PCsrc_MUX(
    input logic PCsrc,
    input logic [31:0] branch_PC,
    input logic [31:0] inc_PC,
    output logic [31:0] next_PC
);




endmodule

