module ImmGen(
    input logic [1:0] ImmSrc,
    input logic [31:0] instruction,
    output logic [31:0] Imm  
);



endmodule
  


